module decoder
#(
	parameter N = 32
)
(
	input      [4:0]  Write_Register_i,
	output reg [N-1:0] Decoder_Out

	
);
	always@(*) begin
	case (Write_Register_i)
	
	0	 : Decoder_Out = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
	1	 : Decoder_Out = 32'b0000_0000_0000_0000_0000_0000_0000_0010;
	2	 : Decoder_Out = 32'b0000_0000_0000_0000_0000_0000_0000_0100;
	3	 : Decoder_Out = 32'b0000_0000_0000_0000_0000_0000_0000_1000;
	4	 : Decoder_Out = 32'b0000_0000_0000_0000_0000_0000_0001_0000;
	5	 : Decoder_Out = 32'b0000_0000_0000_0000_0000_0000_0010_0000;
	6	 : Decoder_Out = 32'b0000_0000_0000_0000_0000_0000_0100_0000;
	7	 : Decoder_Out = 32'b0000_0000_0000_0000_0000_0000_1000_0000;
	8	 : Decoder_Out = 32'b0000_0000_0000_0000_0000_0001_0000_0000;
	9	 : Decoder_Out = 32'b0000_0000_0000_0000_0000_0010_0000_0000;
	10	 : Decoder_Out = 32'b0000_0000_0000_0000_0000_0100_0000_0000;
	11	 : Decoder_Out = 32'b0000_0000_0000_0000_0000_1000_0000_0000;
	12	 : Decoder_Out = 32'b0000_0000_0000_0000_0001_0000_0000_0000;
	13	 : Decoder_Out = 32'b0000_0000_0000_0000_0010_0000_0000_0000;
	14	 : Decoder_Out = 32'b0000_0000_0000_0000_0100_0000_0000_0000;
	15	 : Decoder_Out = 32'b0000_0000_0000_0000_1000_0000_0000_0000;
	16	 : Decoder_Out = 32'b0000_0000_0000_0001_0000_0000_0000_0000;
	17	 : Decoder_Out = 32'b0000_0000_0000_0010_0000_0000_0000_0000;
	18	 : Decoder_Out = 32'b0000_0000_0000_0100_0000_0000_0000_0000;
	19	 : Decoder_Out = 32'b0000_0000_0000_1000_0000_0000_0000_0000;
	20	 : Decoder_Out = 32'b0000_0000_0001_0000_0000_0000_0000_0000;
	21	 : Decoder_Out = 32'b0000_0000_0010_0000_0000_0000_0000_0000;
	22	 : Decoder_Out = 32'b0000_0000_0100_0000_0000_0000_0000_0000;
	23	 : Decoder_Out = 32'b0000_0000_1000_0000_0000_0000_0000_0000;
	24	 : Decoder_Out = 32'b0000_0001_0000_0000_0000_0000_0000_0000;
	25	 : Decoder_Out = 32'b0000_0010_0000_0000_0000_0000_0000_0000;
	26	 : Decoder_Out = 32'b0000_0100_0000_0000_0000_0000_0000_0000;
	27	 : Decoder_Out = 32'b0000_1000_0000_0000_0000_0000_0000_0000;
	28	 : Decoder_Out = 32'b0001_0000_0000_0000_0000_0000_0000_0000;
	29	 : Decoder_Out = 32'b0010_0000_0000_0000_0000_0000_0000_0000;
	30	 : Decoder_Out = 32'b0100_0000_0000_0000_0000_0000_0000_0000;
	31	 : Decoder_Out = 32'b1000_0000_0000_0000_0000_0000_0000_0000;
	

	
	endcase
	end

endmodule 
	
	
	
	

	
	
	
	